//This module controls multi-device acces to synchronous RAM resources

module ramcontroller




endmodule
